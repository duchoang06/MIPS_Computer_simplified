module Exception_Handle
	(
	);
	
endmodule 
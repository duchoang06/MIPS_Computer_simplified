module ALU
	(
		input [3 :0] ALU_control,
		input [31:0] ALU_operand_1,
		input [31:0] ALU_operand_2,
		output [31:0] ALU_result,
		output [7:0] ALU_status
	);
	

	
endmodule 
module ALU_control 
	(
		input [1:0] ALU_control_opcode,
		input [5:0] ALU_control_funct,
		output reg [3:0] ALU_control_out
	);

	always @(ALU_control_opcode, ALU_control_funct) begin
	
	
	
	end
	
endmodule 